module half_adder_tb();
	reg a,b;
	wire s,c;
	initial 


	
